/****************************************************************************
 * uvmdev_delegating_mem.svh
 ****************************************************************************/

/**
 * Class: uvmdev_delegating_mem
 * 
 * Supports delegating memory acceses to one of several memory interfaces
 */
class uvmdev_delegating_mem;

	function new();

	endfunction


endclass


