/****************************************************************************
 * uvmdev_if.svh
 ****************************************************************************/

/**
 * Class: uvmdev_if
 * 
 * TODO: Add class documentation
 */
class uvmdev_if;


endclass


