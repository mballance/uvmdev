/****************************************************************************
 * uvmdev_if.svh
 ****************************************************************************/

/**
 * Class: uvmdev_if
 * 
 * TODO: Add class documentation
 */
interface class uvmdev_if;


endclass


